/*******************************************************************
 *
 * ETF Comment header
 *
 *******************************************************************/

/*******************************************************************
 *
 * Logic gate: NAND -> Y = !(A & B)
 *  
 *     -------------
 *     | A | B | Y |
 *     -------------
 *     | 0 | 0 | 1 |
 *     -------------
 *     | 0 | 1 | 1 |
 *     -------------
 *     | 1 | 0 | 1 |
 *     -------------
 *     | 1 | 1 | 0 |
 *     -------------
 *
 *******************************************************************/
module nand_gate(
    input i_A, 
    input i_B, 
    output o_Y
);
    assign o_Y = ~(i_A & i_B);
    /** Zadatak 1. Ispod unijeti logicku funkciju "NAND" logickog kola! */
    
endmodule

