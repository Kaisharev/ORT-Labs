/*******************************************************************
 *
 * ETF Comment header
 *
 *******************************************************************/

/*******************************************************************
 *
 * Logic gate: NOR -> Y = !(A | B)
 *  
 *     -------------
 *     | A | B | Y |
 *     -------------
 *     | 0 | 0 | 1 |
 *     -------------
 *     | 0 | 1 | 0 |
 *     -------------
 *     | 1 | 0 | 0 |
 *     -------------
 *     | 1 | 1 | 0 |
 *     -------------
 *
 *******************************************************************/
module nor_gate(
    input i_A, 
    input i_B, 
    output o_Y
);
    assign o_Y = ~(i_A | i_B);

    /** Zadatak 3. Ispod unijeti logicku funkciju "NOR" logickog kola! */
    
endmodule

